// Jesus Eduardo Esparza Soto
//Comparador de 4 bits


//Modulo 

module com4b (a,b,res);

		//puertos
		//sentido    tipo  tamaño   nombre
		input              [3:0]    a,b;
		output       reg   [1:0]    res;
		
//Asignaciones


		//secuenciales
		always@(a or b)
		begin 
			if(a>b)
				res=1;
			else if(a<b)
				res=2;
			else
				res=0;
			
		end
endmodule
		